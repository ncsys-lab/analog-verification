* NGSPICE file created from vref_gen_nmos_with_trim.ext - technology: sky130A

.subckt nfet$$185807916 a_4484_n32# a_2832_n32# a_944_n32# li_5147_n4# a_4720_n32#
+ a_n50_0# li_1607_n4# a_6372_n32# li_3023_n4# li_6563_n4# a_6608_n32# li_4439_n4#
+ a_1652_n32# li_427_n4# a_3540_n32# li_5383_n4# a_5192_n32# li_1843_n4# li_6799_n4#
+ li_3259_n4# a_5428_n32# li_663_n4# a_7024_0# a_2360_n32# a_472_n32# li_5619_n4#
+ li_2079_n4# li_3495_n4# a_4248_n32# a_708_n32# a_6136_n32# li_899_n4# a_1180_n32#
+ li_5855_n4# li_2315_n4# li_3731_n4# a_4956_n32# a_3068_n32# a_1416_n32# a_6844_n32#
+ a_3304_n32# li_4675_n4# SUB li_1135_n4# li_2551_n4# li_6091_n4# a_1888_n32# li_3967_n4#
+ a_3776_n32# a_2124_n32# a_5900_n32# a_5664_n32# a_236_n32# a_0_n32# li_4911_n4#
+ a_4012_n32# li_1371_n4# li_2787_n4# li_6327_n4# a_2596_n32# li_191_n4# li_4203_n4#
X0 a_n50_0# a_0_n32# a_n50_0# SUB sky130_fd_pr__nfet_05v0_nvt ad=0.25 pd=2.5 as=25u ps=5m w=1 l=0.4
X1 a_7024_0# a_6844_n32# a_7024_0# SUB sky130_fd_pr__nfet_05v0_nvt ad=0.25 pd=2.5 as=25u ps=5m w=1 l=0.4
.ends

.subckt nfet$$185804844 a_n50_0# a_156_n32# li_111_n4# a_256_0# a_0_n32#
X0 a_n50_0# a_0_n32# a_n50_0# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=2.5 as=25u ps=5m w=1 l=0
X1 a_256_0# a_156_n32# a_256_0# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=2.5 as=25u ps=5m w=1 l=0
.ends

.subckt pfet_symbolic_CDNS_625341251781 a_n50_0# a_0_n26# a_100_0# w_n89_n36#
X0 a_100_0# a_0_n26# a_n50_0# w_n89_n36# sky130_fd_pr__pfet_01v8 ad=0.75 pd=6.5 as=0.75 ps=6.5 w=3 l=0.5
.ends

.subckt pfet_CDNS_625341251780 pfet_symbolic_CDNS_625341251781_0/a_100_0# pfet_symbolic_CDNS_625341251781_0/a_n50_0#
+ w_n119_n66# pfet_symbolic_CDNS_625341251781_0/a_0_n26#
Xpfet_symbolic_CDNS_625341251781_0 pfet_symbolic_CDNS_625341251781_0/a_n50_0# pfet_symbolic_CDNS_625341251781_0/a_0_n26#
+ pfet_symbolic_CDNS_625341251781_0/a_100_0# w_n119_n66# pfet_symbolic_CDNS_625341251781
.ends

.subckt vref_gen_nmos_with_trim trim9 trim10 trim8 trim7 trim6 trim5 trim4 trim3 trim2
+ trim1 vpwr vref vgnd
Xnfet$$185807916_25 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_11728_8706# a_9246_2300# li_11728_8706# vref a_9246_2300# li_11728_8706# a_9246_2300#
+ vref a_9246_2300# li_11728_8706# a_9246_2300# vref li_11728_8706# vref a_9246_2300#
+ li_11728_8706# vref a_9246_2300# a_9246_2300# vref li_11728_8706# li_11728_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_11728_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_11728_8706#
+ li_11728_8706# vref a_9246_2300# li_11728_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_11728_8706# a_9246_2300# vref vref li_11728_8706#
+ a_9246_2300# li_11728_8706# vref nfet$$185807916
Xnfet$$185807916_14 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_8664_8706# a_9246_2300# li_8664_8706# vref a_9246_2300# li_8664_8706# a_9246_2300#
+ vref a_9246_2300# li_8664_8706# a_9246_2300# vref li_8664_8706# vref a_9246_2300#
+ li_8664_8706# vref a_9246_2300# a_9246_2300# vref li_8664_8706# li_8664_8706# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_8664_8706# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_8664_8706# li_8664_8706#
+ vref a_9246_2300# li_8664_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_8664_8706# a_9246_2300# vref vref li_8664_8706# a_9246_2300#
+ li_8664_8706# vref nfet$$185807916
Xnfet$$185804844_2 w_15508_6628# w_15508_7639# w_15508_7639# w_15508_6628# w_15508_7639#
+ nfet$$185804844
Xnfet$$185807916_26 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_13263_8706# a_9246_2300# li_13263_8706# vref a_9246_2300# li_13263_8706# a_9246_2300#
+ vref a_9246_2300# li_13263_8706# a_9246_2300# vref li_13263_8706# vref a_9246_2300#
+ li_13263_8706# vref a_9246_2300# a_9246_2300# vref li_13263_8706# li_13263_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_13263_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_13263_8706#
+ li_13263_8706# vref a_9246_2300# li_13263_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_13263_8706# a_9246_2300# vref vref li_13263_8706#
+ a_9246_2300# li_13263_8706# vref nfet$$185807916
Xnfet$$185807916_15 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_8664_8706# a_9246_2300# li_8664_8706# vref a_9246_2300# li_8664_8706# a_9246_2300#
+ vref a_9246_2300# li_8664_8706# a_9246_2300# vref li_8664_8706# vref a_9246_2300#
+ li_8664_8706# vref a_9246_2300# a_9246_2300# vref li_8664_8706# li_8664_8706# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_8664_8706# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_8664_8706# li_8664_8706#
+ vref a_9246_2300# li_8664_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_8664_8706# a_9246_2300# vref vref li_8664_8706# a_9246_2300#
+ li_8664_8706# vref nfet$$185807916
Xnfet$$185804844_3 w_15508_5617# w_15508_6628# w_15508_6628# w_15508_5617# w_15508_6628#
+ nfet$$185804844
Xnfet$$185807916_27 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_13263_8706# a_9246_2300# li_13263_8706# vref a_9246_2300# li_13263_8706# a_9246_2300#
+ vref a_9246_2300# li_13263_8706# a_9246_2300# vref li_13263_8706# vref a_9246_2300#
+ li_13263_8706# vref a_9246_2300# a_9246_2300# vref li_13263_8706# li_13263_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_13263_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_13263_8706#
+ li_13263_8706# vref a_9246_2300# li_13263_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_13263_8706# a_9246_2300# vref vref li_13263_8706#
+ a_9246_2300# li_13263_8706# vref nfet$$185807916
Xnfet$$185807916_16 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_8664_8706# a_9246_2300# li_8664_8706# vref a_9246_2300# li_8664_8706# a_9246_2300#
+ vref a_9246_2300# li_8664_8706# a_9246_2300# vref li_8664_8706# vref a_9246_2300#
+ li_8664_8706# vref a_9246_2300# a_9246_2300# vref li_8664_8706# li_8664_8706# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_8664_8706# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_8664_8706# li_8664_8706#
+ vref a_9246_2300# li_8664_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_8664_8706# a_9246_2300# vref vref li_8664_8706# a_9246_2300#
+ li_8664_8706# vref nfet$$185807916
Xnfet$$185804844_4 w_15508_2584# w_15508_3595# w_15508_3595# w_15508_2584# w_15508_3595#
+ nfet$$185804844
Xnfet$$185807916_28 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_13263_8706# a_9246_2300# li_13263_8706# vref a_9246_2300# li_13263_8706# a_9246_2300#
+ vref a_9246_2300# li_13263_8706# a_9246_2300# vref li_13263_8706# vref a_9246_2300#
+ li_13263_8706# vref a_9246_2300# a_9246_2300# vref li_13263_8706# li_13263_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_13263_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_13263_8706#
+ li_13263_8706# vref a_9246_2300# li_13263_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_13263_8706# a_9246_2300# vref vref li_13263_8706#
+ a_9246_2300# li_13263_8706# vref nfet$$185807916
Xnfet$$185807916_17 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_8664_8706# a_9246_2300# li_8664_8706# vref a_9246_2300# li_8664_8706# a_9246_2300#
+ vref a_9246_2300# li_8664_8706# a_9246_2300# vref li_8664_8706# vref a_9246_2300#
+ li_8664_8706# vref a_9246_2300# a_9246_2300# vref li_8664_8706# li_8664_8706# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_8664_8706# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_8664_8706# li_8664_8706#
+ vref a_9246_2300# li_8664_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_8664_8706# a_9246_2300# vref vref li_8664_8706# a_9246_2300#
+ li_8664_8706# vref nfet$$185807916
Xnfet$$185804844_5 w_15508_3595# w_15508_4606# w_15508_4606# w_15508_3595# w_15508_4606#
+ nfet$$185804844
Xnfet$$185807916_29 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_13263_8706# a_9246_2300# li_13263_8706# vref a_9246_2300# li_13263_8706# a_9246_2300#
+ vref a_9246_2300# li_13263_8706# a_9246_2300# vref li_13263_8706# vref a_9246_2300#
+ li_13263_8706# vref a_9246_2300# a_9246_2300# vref li_13263_8706# li_13263_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_13263_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_13263_8706#
+ li_13263_8706# vref a_9246_2300# li_13263_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_13263_8706# a_9246_2300# vref vref li_13263_8706#
+ a_9246_2300# li_13263_8706# vref nfet$$185807916
Xnfet$$185807916_18 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_9621_9700# a_9246_2300# li_9621_9700# vref a_9246_2300# li_9621_9700# a_9246_2300#
+ vref a_9246_2300# li_9621_9700# a_9246_2300# vref li_9621_9700# vref a_9246_2300#
+ li_9621_9700# vref a_9246_2300# a_9246_2300# vref li_9621_9700# li_9621_9700# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_9621_9700# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_9621_9700# li_9621_9700#
+ vref a_9246_2300# li_9621_9700# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_9621_9700# a_9246_2300# vref vref li_9621_9700# a_9246_2300#
+ li_9621_9700# vref nfet$$185807916
Xnfet$$185804844_6 w_15508_7639# a_9246_2300# a_9246_2300# w_15508_7639# a_9246_2300#
+ nfet$$185804844
Xnfet$$185807916_19 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_9621_9700# a_9246_2300# li_9621_9700# vref a_9246_2300# li_9621_9700# a_9246_2300#
+ vref a_9246_2300# li_9621_9700# a_9246_2300# vref li_9621_9700# vref a_9246_2300#
+ li_9621_9700# vref a_9246_2300# a_9246_2300# vref li_9621_9700# li_9621_9700# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_9621_9700# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_9621_9700# li_9621_9700#
+ vref a_9246_2300# li_9621_9700# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_9621_9700# a_9246_2300# vref vref li_9621_9700# a_9246_2300#
+ li_9621_9700# vref nfet$$185807916
Xnfet$$185804844_7 w_16618_2584# w_16618_3595# w_16618_3595# w_16618_2584# w_16618_3595#
+ nfet$$185804844
Xnfet$$185804844_8 w_16618_3595# w_16618_4606# w_16618_4606# w_16618_3595# w_16618_4606#
+ nfet$$185804844
Xnfet$$185804844_9 w_16618_4606# w_16618_5617# w_16618_5617# w_16618_4606# w_16618_5617#
+ nfet$$185804844
Xpfet_CDNS_625341251780_0 li_4201_8706# vpwr vpwr trim3 pfet_CDNS_625341251780
Xpfet_CDNS_625341251780_1 li_5606_8706# vpwr vpwr trim4 pfet_CDNS_625341251780
Xpfet_CDNS_625341251780_2 li_3109_8706# vpwr vpwr trim2 pfet_CDNS_625341251780
Xpfet_CDNS_625341251780_3 li_2212_8706# vpwr vpwr trim1 pfet_CDNS_625341251780
Xpfet_CDNS_625341251780_4 li_7153_8706# vpwr vpwr trim5 pfet_CDNS_625341251780
Xpfet_CDNS_625341251780_5 li_8664_8706# vpwr vpwr trim6 pfet_CDNS_625341251780
Xpfet_CDNS_625341251780_6 li_9621_9700# vpwr vpwr trim7 pfet_CDNS_625341251780
Xpfet_CDNS_625341251780_7 li_11728_8706# vpwr vpwr trim8 pfet_CDNS_625341251780
Xpfet_CDNS_625341251780_8 li_13263_8706# vpwr vpwr trim9 pfet_CDNS_625341251780
Xpfet_CDNS_625341251780_9 li_14765_8706# vpwr vpwr trim10 pfet_CDNS_625341251780
Xnfet$$185807916_0 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref li_2212_8706#
+ a_9246_2300# li_2212_8706# vref a_9246_2300# li_2212_8706# a_9246_2300# vref a_9246_2300#
+ li_2212_8706# a_9246_2300# vref li_2212_8706# vref a_9246_2300# li_2212_8706# vref
+ a_9246_2300# a_9246_2300# vref li_2212_8706# li_2212_8706# a_9246_2300# a_9246_2300#
+ a_9246_2300# vref a_9246_2300# li_2212_8706# vref vref a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_2212_8706# li_2212_8706# vref
+ a_9246_2300# li_2212_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# li_2212_8706# a_9246_2300# vref vref li_2212_8706# a_9246_2300# li_2212_8706#
+ vref nfet$$185807916
Xnfet$$185807916_1 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref li_3109_8706#
+ a_9246_2300# li_3109_8706# vref a_9246_2300# li_3109_8706# a_9246_2300# vref a_9246_2300#
+ li_3109_8706# a_9246_2300# vref li_3109_8706# vref a_9246_2300# li_3109_8706# vref
+ a_9246_2300# a_9246_2300# vref li_3109_8706# li_3109_8706# a_9246_2300# a_9246_2300#
+ a_9246_2300# vref a_9246_2300# li_3109_8706# vref vref a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_3109_8706# li_3109_8706# vref
+ a_9246_2300# li_3109_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# li_3109_8706# a_9246_2300# vref vref li_3109_8706# a_9246_2300# li_3109_8706#
+ vref nfet$$185807916
Xnfet$$185807916_2 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref li_3109_8706#
+ a_9246_2300# li_3109_8706# vref a_9246_2300# li_3109_8706# a_9246_2300# vref a_9246_2300#
+ li_3109_8706# a_9246_2300# vref li_3109_8706# vref a_9246_2300# li_3109_8706# vref
+ a_9246_2300# a_9246_2300# vref li_3109_8706# li_3109_8706# a_9246_2300# a_9246_2300#
+ a_9246_2300# vref a_9246_2300# li_3109_8706# vref vref a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_3109_8706# li_3109_8706# vref
+ a_9246_2300# li_3109_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# li_3109_8706# a_9246_2300# vref vref li_3109_8706# a_9246_2300# li_3109_8706#
+ vref nfet$$185807916
Xnfet$$185807916_3 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref li_5606_8706#
+ a_9246_2300# li_5606_8706# vref a_9246_2300# li_5606_8706# a_9246_2300# vref a_9246_2300#
+ li_5606_8706# a_9246_2300# vref li_5606_8706# vref a_9246_2300# li_5606_8706# vref
+ a_9246_2300# a_9246_2300# vref li_5606_8706# li_5606_8706# a_9246_2300# a_9246_2300#
+ a_9246_2300# vref a_9246_2300# li_5606_8706# vref vref a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_5606_8706# li_5606_8706# vref
+ a_9246_2300# li_5606_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# li_5606_8706# a_9246_2300# vref vref li_5606_8706# a_9246_2300# li_5606_8706#
+ vref nfet$$185807916
Xnfet$$185804844_10 w_16618_6628# w_16618_7639# w_16618_7639# w_16618_6628# w_16618_7639#
+ nfet$$185804844
Xnfet$$185807916_4 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref li_5606_8706#
+ a_9246_2300# li_5606_8706# vref a_9246_2300# li_5606_8706# a_9246_2300# vref a_9246_2300#
+ li_5606_8706# a_9246_2300# vref li_5606_8706# vref a_9246_2300# li_5606_8706# vref
+ a_9246_2300# a_9246_2300# vref li_5606_8706# li_5606_8706# a_9246_2300# a_9246_2300#
+ a_9246_2300# vref a_9246_2300# li_5606_8706# vref vref a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_5606_8706# li_5606_8706# vref
+ a_9246_2300# li_5606_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# li_5606_8706# a_9246_2300# vref vref li_5606_8706# a_9246_2300# li_5606_8706#
+ vref nfet$$185807916
Xnfet$$185804844_11 w_16618_5617# w_16618_6628# w_16618_6628# w_16618_5617# w_16618_6628#
+ nfet$$185804844
Xnfet$$185807916_5 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref li_5606_8706#
+ a_9246_2300# li_5606_8706# vref a_9246_2300# li_5606_8706# a_9246_2300# vref a_9246_2300#
+ li_5606_8706# a_9246_2300# vref li_5606_8706# vref a_9246_2300# li_5606_8706# vref
+ a_9246_2300# a_9246_2300# vref li_5606_8706# li_5606_8706# a_9246_2300# a_9246_2300#
+ a_9246_2300# vref a_9246_2300# li_5606_8706# vref vref a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_5606_8706# li_5606_8706# vref
+ a_9246_2300# li_5606_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# li_5606_8706# a_9246_2300# vref vref li_5606_8706# a_9246_2300# li_5606_8706#
+ vref nfet$$185807916
Xnfet$$185804844_12 w_16618_8650# w_15508_2584# w_15508_2584# w_16618_8650# w_15508_2584#
+ nfet$$185804844
Xnfet$$185807916_6 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref li_5606_8706#
+ a_9246_2300# li_5606_8706# vref a_9246_2300# li_5606_8706# a_9246_2300# vref a_9246_2300#
+ li_5606_8706# a_9246_2300# vref li_5606_8706# vref a_9246_2300# li_5606_8706# vref
+ a_9246_2300# a_9246_2300# vref li_5606_8706# li_5606_8706# a_9246_2300# a_9246_2300#
+ a_9246_2300# vref a_9246_2300# li_5606_8706# vref vref a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_5606_8706# li_5606_8706# vref
+ a_9246_2300# li_5606_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# li_5606_8706# a_9246_2300# vref vref li_5606_8706# a_9246_2300# li_5606_8706#
+ vref nfet$$185807916
Xnfet$$185804844_13 w_16618_7639# w_16618_8650# w_16618_8650# w_16618_7639# w_16618_8650#
+ nfet$$185804844
Xnfet$$185807916_7 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref li_4201_8706#
+ a_9246_2300# li_4201_8706# vref a_9246_2300# li_4201_8706# a_9246_2300# vref a_9246_2300#
+ li_4201_8706# a_9246_2300# vref li_4201_8706# vref a_9246_2300# li_4201_8706# vref
+ a_9246_2300# a_9246_2300# vref li_4201_8706# li_4201_8706# a_9246_2300# a_9246_2300#
+ a_9246_2300# vref a_9246_2300# li_4201_8706# vref vref a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_4201_8706# li_4201_8706# vref
+ a_9246_2300# li_4201_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# li_4201_8706# a_9246_2300# vref vref li_4201_8706# a_9246_2300# li_4201_8706#
+ vref nfet$$185807916
Xnfet$$185804844_14 vgnd w_17752_3595# w_17752_3595# vgnd w_17752_3595# nfet$$185804844
Xnfet$$185807916_8 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref li_4201_8706#
+ a_9246_2300# li_4201_8706# vref a_9246_2300# li_4201_8706# a_9246_2300# vref a_9246_2300#
+ li_4201_8706# a_9246_2300# vref li_4201_8706# vref a_9246_2300# li_4201_8706# vref
+ a_9246_2300# a_9246_2300# vref li_4201_8706# li_4201_8706# a_9246_2300# a_9246_2300#
+ a_9246_2300# vref a_9246_2300# li_4201_8706# vref vref a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_4201_8706# li_4201_8706# vref
+ a_9246_2300# li_4201_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# li_4201_8706# a_9246_2300# vref vref li_4201_8706# a_9246_2300# li_4201_8706#
+ vref nfet$$185807916
Xnfet$$185807916_30 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_14765_8706# a_9246_2300# li_14765_8706# vref a_9246_2300# li_14765_8706# a_9246_2300#
+ vref a_9246_2300# li_14765_8706# a_9246_2300# vref li_14765_8706# vref a_9246_2300#
+ li_14765_8706# vref a_9246_2300# a_9246_2300# vref li_14765_8706# li_14765_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_14765_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_14765_8706#
+ li_14765_8706# vref a_9246_2300# li_14765_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_14765_8706# a_9246_2300# vref vref li_14765_8706#
+ a_9246_2300# li_14765_8706# vref nfet$$185807916
Xnfet$$185804844_15 w_17752_3595# w_16618_2584# w_16618_2584# w_17752_3595# w_16618_2584#
+ nfet$$185804844
Xnfet$$185807916_9 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref li_4201_8706#
+ a_9246_2300# li_4201_8706# vref a_9246_2300# li_4201_8706# a_9246_2300# vref a_9246_2300#
+ li_4201_8706# a_9246_2300# vref li_4201_8706# vref a_9246_2300# li_4201_8706# vref
+ a_9246_2300# a_9246_2300# vref li_4201_8706# li_4201_8706# a_9246_2300# a_9246_2300#
+ a_9246_2300# vref a_9246_2300# li_4201_8706# vref vref a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_4201_8706# li_4201_8706# vref
+ a_9246_2300# li_4201_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# li_4201_8706# a_9246_2300# vref vref li_4201_8706# a_9246_2300# li_4201_8706#
+ vref nfet$$185807916
Xnfet$$185807916_31 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_14765_8706# a_9246_2300# li_14765_8706# vref a_9246_2300# li_14765_8706# a_9246_2300#
+ vref a_9246_2300# li_14765_8706# a_9246_2300# vref li_14765_8706# vref a_9246_2300#
+ li_14765_8706# vref a_9246_2300# a_9246_2300# vref li_14765_8706# li_14765_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_14765_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_14765_8706#
+ li_14765_8706# vref a_9246_2300# li_14765_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_14765_8706# a_9246_2300# vref vref li_14765_8706#
+ a_9246_2300# li_14765_8706# vref nfet$$185807916
Xnfet$$185807916_20 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_9621_9700# a_9246_2300# li_9621_9700# vref a_9246_2300# li_9621_9700# a_9246_2300#
+ vref a_9246_2300# li_9621_9700# a_9246_2300# vref li_9621_9700# vref a_9246_2300#
+ li_9621_9700# vref a_9246_2300# a_9246_2300# vref li_9621_9700# li_9621_9700# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_9621_9700# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_9621_9700# li_9621_9700#
+ vref a_9246_2300# li_9621_9700# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_9621_9700# a_9246_2300# vref vref li_9621_9700# a_9246_2300#
+ li_9621_9700# vref nfet$$185807916
Xnfet$$185807916_32 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_14765_8706# a_9246_2300# li_14765_8706# vref a_9246_2300# li_14765_8706# a_9246_2300#
+ vref a_9246_2300# li_14765_8706# a_9246_2300# vref li_14765_8706# vref a_9246_2300#
+ li_14765_8706# vref a_9246_2300# a_9246_2300# vref li_14765_8706# li_14765_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_14765_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_14765_8706#
+ li_14765_8706# vref a_9246_2300# li_14765_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_14765_8706# a_9246_2300# vref vref li_14765_8706#
+ a_9246_2300# li_14765_8706# vref nfet$$185807916
Xnfet$$185807916_21 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_9621_9700# a_9246_2300# li_9621_9700# vref a_9246_2300# li_9621_9700# a_9246_2300#
+ vref a_9246_2300# li_9621_9700# a_9246_2300# vref li_9621_9700# vref a_9246_2300#
+ li_9621_9700# vref a_9246_2300# a_9246_2300# vref li_9621_9700# li_9621_9700# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_9621_9700# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_9621_9700# li_9621_9700#
+ vref a_9246_2300# li_9621_9700# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_9621_9700# a_9246_2300# vref vref li_9621_9700# a_9246_2300#
+ li_9621_9700# vref nfet$$185807916
Xnfet$$185807916_10 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_7153_8706# a_9246_2300# li_7153_8706# vref a_9246_2300# li_7153_8706# a_9246_2300#
+ vref a_9246_2300# li_7153_8706# a_9246_2300# vref li_7153_8706# vref a_9246_2300#
+ li_7153_8706# vref a_9246_2300# a_9246_2300# vref li_7153_8706# li_7153_8706# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_7153_8706# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_7153_8706# li_7153_8706#
+ vref a_9246_2300# li_7153_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_7153_8706# a_9246_2300# vref vref li_7153_8706# a_9246_2300#
+ li_7153_8706# vref nfet$$185807916
Xnfet$$185807916_33 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_14765_8706# a_9246_2300# li_14765_8706# vref a_9246_2300# li_14765_8706# a_9246_2300#
+ vref a_9246_2300# li_14765_8706# a_9246_2300# vref li_14765_8706# vref a_9246_2300#
+ li_14765_8706# vref a_9246_2300# a_9246_2300# vref li_14765_8706# li_14765_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_14765_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_14765_8706#
+ li_14765_8706# vref a_9246_2300# li_14765_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_14765_8706# a_9246_2300# vref vref li_14765_8706#
+ a_9246_2300# li_14765_8706# vref nfet$$185807916
Xnfet$$185807916_22 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_11728_8706# a_9246_2300# li_11728_8706# vref a_9246_2300# li_11728_8706# a_9246_2300#
+ vref a_9246_2300# li_11728_8706# a_9246_2300# vref li_11728_8706# vref a_9246_2300#
+ li_11728_8706# vref a_9246_2300# a_9246_2300# vref li_11728_8706# li_11728_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_11728_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_11728_8706#
+ li_11728_8706# vref a_9246_2300# li_11728_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_11728_8706# a_9246_2300# vref vref li_11728_8706#
+ a_9246_2300# li_11728_8706# vref nfet$$185807916
Xnfet$$185807916_11 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_7153_8706# a_9246_2300# li_7153_8706# vref a_9246_2300# li_7153_8706# a_9246_2300#
+ vref a_9246_2300# li_7153_8706# a_9246_2300# vref li_7153_8706# vref a_9246_2300#
+ li_7153_8706# vref a_9246_2300# a_9246_2300# vref li_7153_8706# li_7153_8706# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_7153_8706# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_7153_8706# li_7153_8706#
+ vref a_9246_2300# li_7153_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_7153_8706# a_9246_2300# vref vref li_7153_8706# a_9246_2300#
+ li_7153_8706# vref nfet$$185807916
Xnfet$$185807916_23 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_11728_8706# a_9246_2300# li_11728_8706# vref a_9246_2300# li_11728_8706# a_9246_2300#
+ vref a_9246_2300# li_11728_8706# a_9246_2300# vref li_11728_8706# vref a_9246_2300#
+ li_11728_8706# vref a_9246_2300# a_9246_2300# vref li_11728_8706# li_11728_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_11728_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_11728_8706#
+ li_11728_8706# vref a_9246_2300# li_11728_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_11728_8706# a_9246_2300# vref vref li_11728_8706#
+ a_9246_2300# li_11728_8706# vref nfet$$185807916
Xnfet$$185807916_12 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_7153_8706# a_9246_2300# li_7153_8706# vref a_9246_2300# li_7153_8706# a_9246_2300#
+ vref a_9246_2300# li_7153_8706# a_9246_2300# vref li_7153_8706# vref a_9246_2300#
+ li_7153_8706# vref a_9246_2300# a_9246_2300# vref li_7153_8706# li_7153_8706# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_7153_8706# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_7153_8706# li_7153_8706#
+ vref a_9246_2300# li_7153_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_7153_8706# a_9246_2300# vref vref li_7153_8706# a_9246_2300#
+ li_7153_8706# vref nfet$$185807916
Xnfet$$185804844_0 a_9246_2300# vref vref a_9246_2300# vref nfet$$185804844
Xnfet$$185807916_24 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_11728_8706# a_9246_2300# li_11728_8706# vref a_9246_2300# li_11728_8706# a_9246_2300#
+ vref a_9246_2300# li_11728_8706# a_9246_2300# vref li_11728_8706# vref a_9246_2300#
+ li_11728_8706# vref a_9246_2300# a_9246_2300# vref li_11728_8706# li_11728_8706#
+ a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# li_11728_8706# vref vref
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_11728_8706#
+ li_11728_8706# vref a_9246_2300# li_11728_8706# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# li_11728_8706# a_9246_2300# vref vref li_11728_8706#
+ a_9246_2300# li_11728_8706# vref nfet$$185807916
Xnfet$$185807916_13 a_9246_2300# a_9246_2300# a_9246_2300# vref a_9246_2300# vref
+ li_7153_8706# a_9246_2300# li_7153_8706# vref a_9246_2300# li_7153_8706# a_9246_2300#
+ vref a_9246_2300# li_7153_8706# a_9246_2300# vref li_7153_8706# vref a_9246_2300#
+ li_7153_8706# vref a_9246_2300# a_9246_2300# vref li_7153_8706# li_7153_8706# a_9246_2300#
+ a_9246_2300# a_9246_2300# vref a_9246_2300# li_7153_8706# vref vref a_9246_2300#
+ a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300# vref vgnd li_7153_8706# li_7153_8706#
+ vref a_9246_2300# li_7153_8706# a_9246_2300# a_9246_2300# a_9246_2300# a_9246_2300#
+ a_9246_2300# a_9246_2300# li_7153_8706# a_9246_2300# vref vref li_7153_8706# a_9246_2300#
+ li_7153_8706# vref nfet$$185807916
Xnfet$$185804844_1 w_15508_4606# w_15508_5617# w_15508_5617# w_15508_4606# w_15508_5617#
+ nfet$$185804844
.ends

