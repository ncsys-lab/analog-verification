

module comparator_latch #
(
  parameter VREF_to_response_time = -1020,
  parameter VREG_to_response_time = -1038,
  parameter const_response_time = 1285,
  parameter VREF_to_tau = 1037,
  parameter VREG_to_tau = -1248,
  parameter const_tau = 1042,
  parameter VREF_to_response_time_lh = -1006,
  parameter VREG_to_response_time_lh = -1752,
  parameter const_response_time_lh = 1185,
  parameter VREF_to_tau_lh = -1115,
  parameter VREG_to_tau_lh = 1131,
  parameter const_tau_lh = 1529
)
(
  input sys_clk,
  input clk,
  input reset,
  input [15-1:0] VREF,
  input [15-1:0] VREG,
  output [39-1:0] out
);

  reg [17-1:0] state_cycle_counter;
  reg [1-1:0] prev_sys_clk;
  reg [39-1:0] o;
  wire [32-1:0] wait_time;
  wire [44-1:0] tau;
  wire [36-1:0] dvdt;
  wire [32-1:0] wait_time_lh;
  wire [46-1:0] tau_lh;
  wire [38-1:0] dodt;
  reg [32-1:0] fsm;
  localparam fsm_init = 0;
  wire [39-1:0] padr_0;
  wire [12-1:0] padr_bits_1;
  assign padr_bits_1 = 0;
  wire [27-1:0] const_2;
  assign const_2 = 55364812;
  assign padr_0 = { const_2, padr_bits_1 };
  assign out = o;
  wire [32-1:0] padl_3;
  wire [3-1:0] padl_bits_4;
  wire [17-1:0] truncR_5;
  wire [96-1:0] truncR_6;
  wire [163-1:0] truncval_7;
  wire [163-1:0] padl_8;
  wire [85-1:0] padl_bits_9;
  wire [85-1:0] padl_10;
  wire [52-1:0] padl_bits_11;
  wire [52-1:0] padr_12;
  wire [2-1:0] padr_bits_13;
  assign padr_bits_13 = 0;
  wire [94-1:0] truncR_14;
  wire [103-1:0] truncval_15;
  wire [103-1:0] padl_16;
  wire [51-1:0] padl_bits_17;
  wire [51-1:0] padr_18;
  wire [36-1:0] padr_bits_19;
  assign padr_bits_19 = 0;
  assign padr_18 = { VREF, padr_bits_19 };
  assign padl_bits_17 = padr_18;
  assign padl_16 = { { 52{ padl_bits_17[50] } }, padl_bits_17 };
  wire [103-1:0] padl_20;
  wire [51-1:0] padl_bits_21;
  wire [51-1:0] padl_22;
  wire [48-1:0] padl_bits_23;
  wire [48-1:0] param_24;
  assign param_24 = VREF_to_response_time;
  assign padl_bits_23 = param_24;
  assign padl_22 = { { 3{ padl_bits_23[47] } }, padl_bits_23 };
  assign padl_bits_21 = padl_22;
  assign padl_20 = { { 52{ padl_bits_21[50] } }, padl_bits_21 };
  assign truncval_15 = padl_16 * padl_20;
  wire [94-1:0] truncval_imm_25;
  assign truncval_imm_25 = { truncval_15[102], truncval_15[92:0] };
  assign truncR_14 = truncval_imm_25;
  wire [50-1:0] truncR_shift_26;
  assign truncR_shift_26 = truncR_14 >>> 44;
  wire [50-1:0] truncR_imm_27;
  assign truncR_imm_27 = (truncR_14[93])? truncR_shift_26[49:0] : truncR_14[93:44];
  assign padr_12 = { truncR_imm_27, padr_bits_13 };
  wire [98-1:0] truncR_28;
  wire [107-1:0] truncval_29;
  wire [107-1:0] padl_30;
  wire [53-1:0] padl_bits_31;
  wire [53-1:0] padr_32;
  wire [38-1:0] padr_bits_33;
  assign padr_bits_33 = 0;
  assign padr_32 = { VREG, padr_bits_33 };
  assign padl_bits_31 = padr_32;
  assign padl_30 = { { 54{ padl_bits_31[52] } }, padl_bits_31 };
  wire [107-1:0] padl_34;
  wire [53-1:0] padl_bits_35;
  wire [53-1:0] padl_36;
  wire [50-1:0] padl_bits_37;
  wire [50-1:0] param_38;
  assign param_38 = VREG_to_response_time;
  assign padl_bits_37 = param_38;
  assign padl_36 = { { 3{ padl_bits_37[49] } }, padl_bits_37 };
  assign padl_bits_35 = padl_36;
  assign padl_34 = { { 54{ padl_bits_35[52] } }, padl_bits_35 };
  assign truncval_29 = padl_30 * padl_34;
  wire [98-1:0] truncval_imm_39;
  assign truncval_imm_39 = { truncval_29[106], truncval_29[96:0] };
  assign truncR_28 = truncval_imm_39;
  wire [52-1:0] truncR_shift_40;
  assign truncR_shift_40 = truncR_28 >>> 46;
  wire [52-1:0] truncR_imm_41;
  assign truncR_imm_41 = (truncR_28[97])? truncR_shift_40[51:0] : truncR_28[97:46];
  wire [52-1:0] padr_42;
  wire [8-1:0] padr_bits_43;
  assign padr_bits_43 = 0;
  wire [44-1:0] padl_44;
  wire [43-1:0] padl_bits_45;
  wire [1-1:0] toSInt_46;
  assign toSInt_46 = 0;
  wire [43-1:0] toSInt_imm_47;
  wire [42-1:0] param_48;
  assign param_48 = const_response_time;
  assign toSInt_imm_47 = { toSInt_46, param_48 };
  assign padl_bits_45 = toSInt_imm_47;
  assign padl_44 = { { 1{ padl_bits_45[42] } }, padl_bits_45 };
  assign padr_42 = { padl_44, padr_bits_43 };
  assign padl_bits_11 = padr_12 + truncR_imm_41 + padr_42;
  assign padl_10 = { { 33{ padl_bits_11[51] } }, padl_bits_11 };
  assign padl_bits_9 = padl_10;
  assign padl_8 = { { 78{ padl_bits_9[84] } }, padl_bits_9 };
  wire [163-1:0] padl_49;
  wire [85-1:0] padl_bits_50;
  wire [85-1:0] padr_51;
  wire [50-1:0] padr_bits_52;
  assign padr_bits_52 = 0;
  wire [1-1:0] toSInt_53;
  assign toSInt_53 = 0;
  wire [35-1:0] toSInt_imm_54;
  wire [34-1:0] const_55;
  assign const_55 = 78125000;
  assign toSInt_imm_54 = { toSInt_53, const_55 };
  assign padr_51 = { toSInt_imm_54, padr_bits_52 };
  assign padl_bits_50 = padr_51;
  assign padl_49 = { { 78{ padl_bits_50[84] } }, padl_bits_50 };
  assign truncval_7 = padl_8 * padl_49;
  assign truncR_6 = truncval_7[95:0];
  assign truncR_5 = truncR_6[95:79];
  assign padl_bits_4 = truncR_5[16:14];
  wire [29-1:0] padl_bits_zero_56;
  assign padl_bits_zero_56 = 0;
  assign padl_3 = { padl_bits_zero_56, padl_bits_4 };
  assign wait_time = padl_3;
  wire [39-1:0] padr_57;
  wire [12-1:0] padr_bits_58;
  assign padr_bits_58 = 0;
  wire [27-1:0] const_59;
  assign const_59 = 55364812;
  assign padr_57 = { const_59, padr_bits_58 };
  wire [45-1:0] truncR_60;
  wire [46-1:0] truncval_61;
  wire [47-1:0] toUsInt_62;
  wire [88-1:0] truncR_63;
  wire [97-1:0] truncval_64;
  wire [97-1:0] padl_65;
  wire [48-1:0] padl_bits_66;
  wire [48-1:0] padr_67;
  wire [33-1:0] padr_bits_68;
  assign padr_bits_68 = 0;
  assign padr_67 = { VREF, padr_bits_68 };
  assign padl_bits_66 = padr_67;
  assign padl_65 = { { 49{ padl_bits_66[47] } }, padl_bits_66 };
  wire [97-1:0] padl_69;
  wire [48-1:0] padl_bits_70;
  wire [48-1:0] padl_71;
  wire [44-1:0] padl_bits_72;
  wire [1-1:0] toSInt_73;
  assign toSInt_73 = 0;
  wire [44-1:0] toSInt_imm_74;
  wire [43-1:0] param_75;
  assign param_75 = VREF_to_tau;
  assign toSInt_imm_74 = { toSInt_73, param_75 };
  assign padl_bits_72 = toSInt_imm_74;
  assign padl_71 = { { 4{ padl_bits_72[43] } }, padl_bits_72 };
  assign padl_bits_70 = padl_71;
  assign padl_69 = { { 49{ padl_bits_70[47] } }, padl_bits_70 };
  assign truncval_64 = padl_65 * padl_69;
  wire [88-1:0] truncval_imm_76;
  assign truncval_imm_76 = { truncval_64[96], truncval_64[86:0] };
  assign truncR_63 = truncval_imm_76;
  wire [47-1:0] truncR_shift_77;
  assign truncR_shift_77 = truncR_63 >>> 41;
  wire [47-1:0] truncR_imm_78;
  assign truncR_imm_78 = (truncR_63[87])? truncR_shift_77[46:0] : truncR_63[87:41];
  wire [47-1:0] padr_79;
  wire [1-1:0] padr_bits_80;
  assign padr_bits_80 = 0;
  wire [88-1:0] truncR_81;
  wire [97-1:0] truncval_82;
  wire [97-1:0] padl_83;
  wire [48-1:0] padl_bits_84;
  wire [48-1:0] padr_85;
  wire [33-1:0] padr_bits_86;
  assign padr_bits_86 = 0;
  assign padr_85 = { VREG, padr_bits_86 };
  assign padl_bits_84 = padr_85;
  assign padl_83 = { { 49{ padl_bits_84[47] } }, padl_bits_84 };
  wire [97-1:0] padl_87;
  wire [48-1:0] padl_bits_88;
  wire [48-1:0] padl_89;
  wire [45-1:0] padl_bits_90;
  wire [45-1:0] param_91;
  assign param_91 = VREG_to_tau;
  assign padl_bits_90 = param_91;
  assign padl_89 = { { 3{ padl_bits_90[44] } }, padl_bits_90 };
  assign padl_bits_88 = padl_89;
  assign padl_87 = { { 49{ padl_bits_88[47] } }, padl_bits_88 };
  assign truncval_82 = padl_83 * padl_87;
  wire [88-1:0] truncval_imm_92;
  assign truncval_imm_92 = { truncval_82[96], truncval_82[86:0] };
  assign truncR_81 = truncval_imm_92;
  wire [46-1:0] truncR_shift_93;
  assign truncR_shift_93 = truncR_81 >>> 42;
  wire [46-1:0] truncR_imm_94;
  assign truncR_imm_94 = (truncR_81[87])? truncR_shift_93[45:0] : truncR_81[87:42];
  assign padr_79 = { truncR_imm_94, padr_bits_80 };
  wire [47-1:0] padr_95;
  wire [4-1:0] padr_bits_96;
  assign padr_bits_96 = 0;
  wire [43-1:0] padl_97;
  wire [42-1:0] padl_bits_98;
  wire [1-1:0] toSInt_99;
  assign toSInt_99 = 0;
  wire [42-1:0] toSInt_imm_100;
  wire [41-1:0] param_101;
  assign param_101 = const_tau;
  assign toSInt_imm_100 = { toSInt_99, param_101 };
  assign padl_bits_98 = toSInt_imm_100;
  assign padl_97 = { { 1{ padl_bits_98[41] } }, padl_bits_98 };
  assign padr_95 = { padl_97, padr_bits_96 };
  assign toUsInt_62 = truncR_imm_78 + padr_79 + padr_95;
  assign truncval_61 = toUsInt_62[43:0];
  assign truncR_60 = truncval_61[44:0];
  assign tau = truncR_60[44:1];
  wire [39-1:0] padr_102;
  wire [24-1:0] padr_bits_103;
  assign padr_bits_103 = 0;
  wire [16-1:0] toUsInt_104;
  wire [16-1:0] padr_105;
  wire [5-1:0] padr_bits_106;
  assign padr_bits_106 = 0;
  wire [12-1:0] truncval_107;
  wire [12-1:0] padl_108;
  wire [11-1:0] padl_bits_109;
  wire [40-1:0] truncR_110;
  wire [1-1:0] toSInt_111;
  assign toSInt_111 = 0;
  wire [40-1:0] toSInt_imm_112;
  assign toSInt_imm_112 = { toSInt_111, o };
  assign truncR_110 = toSInt_imm_112;
  wire [11-1:0] truncR_shift_113;
  assign truncR_shift_113 = truncR_110 >>> 29;
  wire [11-1:0] truncR_imm_114;
  assign truncR_imm_114 = (truncR_110[39])? truncR_shift_113[10:0] : truncR_110[39:29];
  assign padl_bits_109 = truncR_imm_114;
  assign padl_108 = { { 1{ padl_bits_109[10] } }, padl_bits_109 };
  assign truncval_107 = padl_108;
  wire [11-1:0] truncval_imm_115;
  assign truncval_imm_115 = { truncval_107[11], truncval_107[9:0] };
  assign padr_105 = { truncval_imm_115, padr_bits_106 };
  assign toUsInt_104 = padr_105;
  assign padr_102 = { toUsInt_104[12:0], padr_bits_103 };
  wire [36-1:0] padl_116;
  wire [16-1:0] padl_bits_117;
  wire [36-1:0] truncR_118;
  wire [60-1:0] truncR_119;
  wire [93-1:0] truncval_120;
  wire [93-1:0] padl_121;
  wire [46-1:0] padl_bits_122;
  wire [46-1:0] padl_123;
  wire [16-1:0] padl_bits_124;
  wire [16-1:0] neg_imm_125;
  wire [16-1:0] padr_126;
  wire [5-1:0] padr_bits_127;
  assign padr_bits_127 = 0;
  wire [12-1:0] truncval_128;
  wire [12-1:0] padl_129;
  wire [11-1:0] padl_bits_130;
  wire [40-1:0] truncR_131;
  wire [1-1:0] toSInt_132;
  assign toSInt_132 = 0;
  wire [40-1:0] toSInt_imm_133;
  assign toSInt_imm_133 = { toSInt_132, o };
  assign truncR_131 = toSInt_imm_133;
  wire [11-1:0] truncR_shift_134;
  assign truncR_shift_134 = truncR_131 >>> 29;
  wire [11-1:0] truncR_imm_135;
  assign truncR_imm_135 = (truncR_131[39])? truncR_shift_134[10:0] : truncR_131[39:29];
  assign padl_bits_130 = truncR_imm_135;
  assign padl_129 = { { 1{ padl_bits_130[10] } }, padl_bits_130 };
  assign truncval_128 = padl_129;
  wire [11-1:0] truncval_imm_136;
  assign truncval_imm_136 = { truncval_128[11], truncval_128[9:0] };
  assign padr_126 = { truncval_imm_136, padr_bits_127 };
  assign neg_imm_125 = -padr_126;
  assign padl_bits_124 = neg_imm_125;
  assign padl_123 = { { 30{ padl_bits_124[15] } }, padl_bits_124 };
  assign padl_bits_122 = padl_123;
  assign padl_121 = { { 47{ padl_bits_122[45] } }, padl_bits_122 };
  wire [93-1:0] padl_137;
  wire [46-1:0] padl_bits_138;
  wire [46-1:0] padr_139;
  wire [12-1:0] padr_bits_140;
  assign padr_bits_140 = 0;
  wire [1-1:0] toSInt_141;
  assign toSInt_141 = 0;
  wire [34-1:0] toSInt_imm_142;
  wire [44-1:0] truncval_143;
  assign truncval_143 = 45'd17592186044416 / tau;
  assign toSInt_imm_142 = { toSInt_141, truncval_143[32:0] };
  assign padr_139 = { toSInt_imm_142, padr_bits_140 };
  assign padl_bits_138 = padr_139;
  assign padl_137 = { { 47{ padl_bits_138[45] } }, padl_bits_138 };
  assign truncval_120 = padl_121 * padl_137;
  wire [60-1:0] truncval_imm_144;
  assign truncval_imm_144 = { truncval_120[92], truncval_120[58:0] };
  assign truncR_119 = truncval_imm_144;
  wire [36-1:0] truncR_shift_145;
  assign truncR_shift_145 = truncR_119 >>> 24;
  wire [36-1:0] truncR_imm_146;
  assign truncR_imm_146 = (truncR_119[59])? truncR_shift_145[35:0] : truncR_119[59:24];
  assign truncR_118 = truncR_imm_146;
  wire [16-1:0] truncR_shift_147;
  assign truncR_shift_147 = truncR_118 >>> 20;
  wire [16-1:0] truncR_imm_148;
  assign truncR_imm_148 = (truncR_118[35])? truncR_shift_147[15:0] : truncR_118[35:20];
  assign padl_bits_117 = truncR_imm_148;
  assign padl_116 = { { 20{ padl_bits_117[15] } }, padl_bits_117 };
  assign dvdt = padl_116;
  wire [41-1:0] truncval_149;
  wire [41-1:0] padr_150;
  wire [29-1:0] padr_bits_151;
  assign padr_bits_151 = 0;
  wire [19-1:0] truncR_152;
  wire [19-1:0] padl_153;
  wire [16-1:0] padl_bits_154;
  wire [100-1:0] truncR_155;
  wire [171-1:0] truncval_156;
  wire [171-1:0] padl_157;
  wire [95-1:0] padl_bits_158;
  wire [95-1:0] padl_159;
  wire [60-1:0] padl_bits_160;
  wire [1-1:0] toSInt_161;
  assign toSInt_161 = 0;
  wire [60-1:0] toSInt_imm_162;
  wire [59-1:0] const_163;
  assign const_163 = 57646075;
  assign toSInt_imm_162 = { toSInt_161, const_163 };
  assign padl_bits_160 = toSInt_imm_162;
  assign padl_159 = { { 35{ padl_bits_160[59] } }, padl_bits_160 };
  assign padl_bits_158 = padl_159;
  assign padl_157 = { { 76{ padl_bits_158[94] } }, padl_bits_158 };
  wire [171-1:0] padl_164;
  wire [95-1:0] padl_bits_165;
  wire [95-1:0] padr_166;
  wire [59-1:0] padr_bits_167;
  assign padr_bits_167 = 0;
  assign padr_166 = { dvdt, padr_bits_167 };
  assign padl_bits_165 = padr_166;
  assign padl_164 = { { 76{ padl_bits_165[94] } }, padl_bits_165 };
  assign truncval_156 = padl_157 * padl_164;
  wire [100-1:0] truncval_imm_168;
  assign truncval_imm_168 = { truncval_156[170], truncval_156[98:0] };
  assign truncR_155 = truncval_imm_168;
  wire [16-1:0] truncR_shift_169;
  assign truncR_shift_169 = truncR_155 >>> 84;
  wire [16-1:0] truncR_imm_170;
  assign truncR_imm_170 = (truncR_155[99])? truncR_shift_169[15:0] : truncR_155[99:84];
  assign padl_bits_154 = truncR_imm_170;
  assign padl_153 = { { 3{ padl_bits_154[15] } }, padl_bits_154 };
  assign truncR_152 = padl_153;
  wire [12-1:0] truncR_shift_171;
  assign truncR_shift_171 = truncR_152 >>> 7;
  wire [12-1:0] truncR_imm_172;
  assign truncR_imm_172 = (truncR_152[18])? truncR_shift_171[11:0] : truncR_152[18:7];
  assign padr_150 = { truncR_imm_172, padr_bits_151 };
  assign truncval_149 = padr_150;
  wire [39-1:0] truncval_imm_173;
  assign truncval_imm_173 = { truncval_149[40], truncval_149[37:0] };
  wire [32-1:0] padl_174;
  wire [2-1:0] padl_bits_175;
  wire [16-1:0] truncR_176;
  wire [93-1:0] truncR_177;
  wire [161-1:0] truncval_178;
  wire [161-1:0] padl_179;
  wire [84-1:0] padl_bits_180;
  wire [84-1:0] padl_181;
  wire [51-1:0] padl_bits_182;
  wire [51-1:0] padr_183;
  wire [1-1:0] padr_bits_184;
  assign padr_bits_184 = 0;
  wire [94-1:0] truncR_185;
  wire [103-1:0] truncval_186;
  wire [103-1:0] padl_187;
  wire [51-1:0] padl_bits_188;
  wire [51-1:0] padr_189;
  wire [39-1:0] padr_bits_190;
  assign padr_bits_190 = 0;
  wire [15-1:0] truncR_191;
  assign truncR_191 = VREF;
  wire [12-1:0] truncR_shift_192;
  assign truncR_shift_192 = truncR_191 >>> 3;
  wire [12-1:0] truncR_imm_193;
  assign truncR_imm_193 = (truncR_191[14])? truncR_shift_192[11:0] : truncR_191[14:3];
  assign padr_189 = { truncR_imm_193, padr_bits_190 };
  assign padl_bits_188 = padr_189;
  assign padl_187 = { { 52{ padl_bits_188[50] } }, padl_bits_188 };
  wire [103-1:0] padl_194;
  wire [51-1:0] padl_bits_195;
  wire [51-1:0] padl_196;
  wire [48-1:0] padl_bits_197;
  wire [48-1:0] param_198;
  assign param_198 = VREF_to_response_time_lh;
  assign padl_bits_197 = param_198;
  assign padl_196 = { { 3{ padl_bits_197[47] } }, padl_bits_197 };
  assign padl_bits_195 = padl_196;
  assign padl_194 = { { 52{ padl_bits_195[50] } }, padl_bits_195 };
  assign truncval_186 = padl_187 * padl_194;
  wire [94-1:0] truncval_imm_199;
  assign truncval_imm_199 = { truncval_186[102], truncval_186[92:0] };
  assign truncR_185 = truncval_imm_199;
  wire [50-1:0] truncR_shift_200;
  assign truncR_shift_200 = truncR_185 >>> 44;
  wire [50-1:0] truncR_imm_201;
  assign truncR_imm_201 = (truncR_185[93])? truncR_shift_200[49:0] : truncR_185[93:44];
  assign padr_183 = { truncR_imm_201, padr_bits_184 };
  wire [98-1:0] truncR_202;
  wire [107-1:0] truncval_203;
  wire [107-1:0] padl_204;
  wire [53-1:0] padl_bits_205;
  wire [53-1:0] padr_206;
  wire [41-1:0] padr_bits_207;
  assign padr_bits_207 = 0;
  assign padr_206 = { VREG, padr_bits_207 };
  assign padl_bits_205 = padr_206;
  assign padl_204 = { { 54{ padl_bits_205[52] } }, padl_bits_205 };
  wire [107-1:0] padl_208;
  wire [53-1:0] padl_bits_209;
  wire [53-1:0] padl_210;
  wire [50-1:0] padl_bits_211;
  wire [50-1:0] param_212;
  assign param_212 = VREG_to_response_time_lh;
  assign padl_bits_211 = param_212;
  assign padl_210 = { { 3{ padl_bits_211[49] } }, padl_bits_211 };
  assign padl_bits_209 = padl_210;
  assign padl_208 = { { 54{ padl_bits_209[52] } }, padl_bits_209 };
  assign truncval_203 = padl_204 * padl_208;
  wire [98-1:0] truncval_imm_213;
  assign truncval_imm_213 = { truncval_203[106], truncval_203[96:0] };
  assign truncR_202 = truncval_imm_213;
  wire [51-1:0] truncR_shift_214;
  assign truncR_shift_214 = truncR_202 >>> 47;
  wire [51-1:0] truncR_imm_215;
  assign truncR_imm_215 = (truncR_202[97])? truncR_shift_214[50:0] : truncR_202[97:47];
  wire [51-1:0] padr_216;
  wire [6-1:0] padr_bits_217;
  assign padr_bits_217 = 0;
  wire [45-1:0] padl_218;
  wire [44-1:0] padl_bits_219;
  wire [1-1:0] toSInt_220;
  assign toSInt_220 = 0;
  wire [44-1:0] toSInt_imm_221;
  wire [43-1:0] param_222;
  assign param_222 = const_response_time_lh;
  assign toSInt_imm_221 = { toSInt_220, param_222 };
  assign padl_bits_219 = toSInt_imm_221;
  assign padl_218 = { { 1{ padl_bits_219[43] } }, padl_bits_219 };
  assign padr_216 = { padl_218, padr_bits_217 };
  assign padl_bits_182 = padr_183 + truncR_imm_215 + padr_216;
  assign padl_181 = { { 33{ padl_bits_182[50] } }, padl_bits_182 };
  assign padl_bits_180 = padl_181;
  assign padl_179 = { { 77{ padl_bits_180[83] } }, padl_bits_180 };
  wire [161-1:0] padl_223;
  wire [84-1:0] padl_bits_224;
  wire [84-1:0] padr_225;
  wire [49-1:0] padr_bits_226;
  assign padr_bits_226 = 0;
  wire [1-1:0] toSInt_227;
  assign toSInt_227 = 0;
  wire [35-1:0] toSInt_imm_228;
  wire [34-1:0] const_229;
  assign const_229 = 78125000;
  assign toSInt_imm_228 = { toSInt_227, const_229 };
  assign padr_225 = { toSInt_imm_228, padr_bits_226 };
  assign padl_bits_224 = padr_225;
  assign padl_223 = { { 77{ padl_bits_224[83] } }, padl_bits_224 };
  assign truncval_178 = padl_179 * padl_223;
  assign truncR_177 = truncval_178[92:0];
  assign truncR_176 = truncR_177[92:77];
  assign padl_bits_175 = truncR_176[15:14];
  wire [30-1:0] padl_bits_zero_230;
  assign padl_bits_zero_230 = 0;
  assign padl_174 = { padl_bits_zero_230, padl_bits_175 };
  assign wait_time_lh = padl_174;
  wire [39-1:0] padl_231;
  wire [36-1:0] padl_bits_232;
  wire [36-1:0] const_233;
  assign const_233 = 68719476;
  assign padl_bits_232 = const_233;
  wire [3-1:0] padl_bits_zero_234;
  assign padl_bits_zero_234 = 0;
  assign padl_231 = { padl_bits_zero_234, padl_bits_232 };
  wire [49-1:0] truncR_235;
  wire [50-1:0] truncval_236;
  wire [51-1:0] toUsInt_237;
  wire [96-1:0] truncR_238;
  wire [105-1:0] truncval_239;
  wire [105-1:0] padl_240;
  wire [52-1:0] padl_bits_241;
  wire [52-1:0] padr_242;
  wire [40-1:0] padr_bits_243;
  assign padr_bits_243 = 0;
  wire [15-1:0] truncR_244;
  assign truncR_244 = VREF;
  wire [12-1:0] truncR_shift_245;
  assign truncR_shift_245 = truncR_244 >>> 3;
  wire [12-1:0] truncR_imm_246;
  assign truncR_imm_246 = (truncR_244[14])? truncR_shift_245[11:0] : truncR_244[14:3];
  assign padr_242 = { truncR_imm_246, padr_bits_243 };
  assign padl_bits_241 = padr_242;
  assign padl_240 = { { 53{ padl_bits_241[51] } }, padl_bits_241 };
  wire [105-1:0] padl_247;
  wire [52-1:0] padl_bits_248;
  wire [52-1:0] padl_249;
  wire [49-1:0] padl_bits_250;
  wire [49-1:0] param_251;
  assign param_251 = VREF_to_tau_lh;
  assign padl_bits_250 = param_251;
  assign padl_249 = { { 3{ padl_bits_250[48] } }, padl_bits_250 };
  assign padl_bits_248 = padl_249;
  assign padl_247 = { { 53{ padl_bits_248[51] } }, padl_bits_248 };
  assign truncval_239 = padl_240 * padl_247;
  wire [96-1:0] truncval_imm_252;
  assign truncval_imm_252 = { truncval_239[104], truncval_239[94:0] };
  assign truncR_238 = truncval_imm_252;
  wire [51-1:0] truncR_shift_253;
  assign truncR_shift_253 = truncR_238 >>> 45;
  wire [51-1:0] truncR_imm_254;
  assign truncR_imm_254 = (truncR_238[95])? truncR_shift_253[50:0] : truncR_238[95:45];
  wire [51-1:0] padr_255;
  wire [3-1:0] padr_bits_256;
  assign padr_bits_256 = 0;
  wire [90-1:0] truncR_257;
  wire [99-1:0] truncval_258;
  wire [99-1:0] padl_259;
  wire [49-1:0] padl_bits_260;
  wire [49-1:0] padr_261;
  wire [37-1:0] padr_bits_262;
  assign padr_bits_262 = 0;
  assign padr_261 = { VREG, padr_bits_262 };
  assign padl_bits_260 = padr_261;
  assign padl_259 = { { 50{ padl_bits_260[48] } }, padl_bits_260 };
  wire [99-1:0] padl_263;
  wire [49-1:0] padl_bits_264;
  wire [49-1:0] padl_265;
  wire [45-1:0] padl_bits_266;
  wire [1-1:0] toSInt_267;
  assign toSInt_267 = 0;
  wire [45-1:0] toSInt_imm_268;
  wire [44-1:0] param_269;
  assign param_269 = VREG_to_tau_lh;
  assign toSInt_imm_268 = { toSInt_267, param_269 };
  assign padl_bits_266 = toSInt_imm_268;
  assign padl_265 = { { 4{ padl_bits_266[44] } }, padl_bits_266 };
  assign padl_bits_264 = padl_265;
  assign padl_263 = { { 50{ padl_bits_264[48] } }, padl_bits_264 };
  assign truncval_258 = padl_259 * padl_263;
  wire [90-1:0] truncval_imm_270;
  assign truncval_imm_270 = { truncval_258[98], truncval_258[88:0] };
  assign truncR_257 = truncval_imm_270;
  wire [48-1:0] truncR_shift_271;
  assign truncR_shift_271 = truncR_257 >>> 42;
  wire [48-1:0] truncR_imm_272;
  assign truncR_imm_272 = (truncR_257[89])? truncR_shift_271[47:0] : truncR_257[89:42];
  assign padr_255 = { truncR_imm_272, padr_bits_256 };
  wire [51-1:0] padr_273;
  wire [6-1:0] padr_bits_274;
  assign padr_bits_274 = 0;
  wire [45-1:0] padl_275;
  wire [44-1:0] padl_bits_276;
  wire [1-1:0] toSInt_277;
  assign toSInt_277 = 0;
  wire [44-1:0] toSInt_imm_278;
  wire [43-1:0] param_279;
  assign param_279 = const_tau_lh;
  assign toSInt_imm_278 = { toSInt_277, param_279 };
  assign padl_bits_276 = toSInt_imm_278;
  assign padl_275 = { { 1{ padl_bits_276[43] } }, padl_bits_276 };
  assign padr_273 = { padl_275, padr_bits_274 };
  assign toUsInt_237 = truncR_imm_254 + padr_255 + padr_273;
  assign truncval_236 = toUsInt_237[47:0];
  assign truncR_235 = truncval_236[48:0];
  assign tau_lh = truncR_235[48:3];
  wire [39-1:0] padr_280;
  wire [24-1:0] padr_bits_281;
  assign padr_bits_281 = 0;
  wire [16-1:0] toUsInt_282;
  wire [34-1:0] truncR_283;
  wire [35-1:0] truncval_284;
  wire [35-1:0] padl_285;
  wire [34-1:0] padl_bits_286;
  wire [40-1:0] truncR_287;
  wire [1-1:0] toSInt_288;
  assign toSInt_288 = 0;
  wire [40-1:0] toSInt_imm_289;
  assign toSInt_imm_289 = { toSInt_288, o };
  assign truncR_287 = toSInt_imm_289;
  wire [34-1:0] truncR_shift_290;
  assign truncR_shift_290 = truncR_287 >>> 6;
  wire [34-1:0] truncR_imm_291;
  assign truncR_imm_291 = (truncR_287[39])? truncR_shift_290[33:0] : truncR_287[39:6];
  assign padl_bits_286 = truncR_imm_291;
  assign padl_285 = { { 1{ padl_bits_286[33] } }, padl_bits_286 };
  assign truncval_284 = padl_285;
  wire [34-1:0] truncval_imm_292;
  assign truncval_imm_292 = { truncval_284[34], truncval_284[32:0] };
  assign truncR_283 = truncval_imm_292;
  wire [16-1:0] truncR_shift_293;
  assign truncR_shift_293 = truncR_283 >>> 18;
  wire [16-1:0] truncR_imm_294;
  assign truncR_imm_294 = (truncR_283[33])? truncR_shift_293[15:0] : truncR_283[33:18];
  assign toUsInt_282 = truncR_imm_294;
  assign padr_280 = { toUsInt_282[12:0], padr_bits_281 };
  wire [38-1:0] padl_295;
  wire [17-1:0] padl_bits_296;
  wire [38-1:0] truncR_297;
  wire [98-1:0] truncR_298;
  wire [129-1:0] truncval_299;
  wire [129-1:0] padl_300;
  wire [64-1:0] padl_bits_301;
  wire [64-1:0] padl_302;
  wire [35-1:0] padl_bits_303;
  wire [35-1:0] padr_304;
  wire [6-1:0] padr_bits_305;
  assign padr_bits_305 = 0;
  wire [29-1:0] padl_306;
  wire [28-1:0] padl_bits_307;
  wire [1-1:0] toSInt_308;
  assign toSInt_308 = 0;
  wire [28-1:0] toSInt_imm_309;
  wire [27-1:0] const_310;
  assign const_310 = 55364812;
  assign toSInt_imm_309 = { toSInt_308, const_310 };
  assign padl_bits_307 = toSInt_imm_309;
  assign padl_306 = { { 1{ padl_bits_307[27] } }, padl_bits_307 };
  assign padr_304 = { padl_306, padr_bits_305 };
  wire [35-1:0] padl_311;
  wire [34-1:0] padl_bits_312;
  wire [40-1:0] truncR_313;
  wire [1-1:0] toSInt_314;
  assign toSInt_314 = 0;
  wire [40-1:0] toSInt_imm_315;
  assign toSInt_imm_315 = { toSInt_314, o };
  assign truncR_313 = toSInt_imm_315;
  wire [34-1:0] truncR_shift_316;
  assign truncR_shift_316 = truncR_313 >>> 6;
  wire [34-1:0] truncR_imm_317;
  assign truncR_imm_317 = (truncR_313[39])? truncR_shift_316[33:0] : truncR_313[39:6];
  assign padl_bits_312 = truncR_imm_317;
  assign padl_311 = { { 1{ padl_bits_312[33] } }, padl_bits_312 };
  assign padl_bits_303 = padr_304 - padl_311;
  assign padl_302 = { { 29{ padl_bits_303[34] } }, padl_bits_303 };
  assign padl_bits_301 = padl_302;
  assign padl_300 = { { 65{ padl_bits_301[63] } }, padl_bits_301 };
  wire [129-1:0] padl_318;
  wire [64-1:0] padl_bits_319;
  wire [64-1:0] padr_320;
  wire [30-1:0] padr_bits_321;
  assign padr_bits_321 = 0;
  wire [1-1:0] toSInt_322;
  assign toSInt_322 = 0;
  wire [34-1:0] toSInt_imm_323;
  wire [46-1:0] truncval_324;
  assign truncval_324 = 47'd70368744177664 / tau_lh;
  assign toSInt_imm_323 = { toSInt_322, truncval_324[32:0] };
  assign padr_320 = { toSInt_imm_323, padr_bits_321 };
  assign padl_bits_319 = padr_320;
  assign padl_318 = { { 65{ padl_bits_319[63] } }, padl_bits_319 };
  assign truncval_299 = padl_300 * padl_318;
  wire [98-1:0] truncval_imm_325;
  assign truncval_imm_325 = { truncval_299[128], truncval_299[96:0] };
  assign truncR_298 = truncval_imm_325;
  wire [38-1:0] truncR_shift_326;
  assign truncR_shift_326 = truncR_298 >>> 60;
  wire [38-1:0] truncR_imm_327;
  assign truncR_imm_327 = (truncR_298[97])? truncR_shift_326[37:0] : truncR_298[97:60];
  assign truncR_297 = truncR_imm_327;
  wire [17-1:0] truncR_shift_328;
  assign truncR_shift_328 = truncR_297 >>> 21;
  wire [17-1:0] truncR_imm_329;
  assign truncR_imm_329 = (truncR_297[37])? truncR_shift_328[16:0] : truncR_297[37:21];
  assign padl_bits_296 = truncR_imm_329;
  assign padl_295 = { { 21{ padl_bits_296[16] } }, padl_bits_296 };
  assign dodt = padl_295;
  wire [41-1:0] truncval_330;
  wire [41-1:0] padr_331;
  wire [6-1:0] padr_bits_332;
  assign padr_bits_332 = 0;
  wire [35-1:0] padr_333;
  wire [17-1:0] padr_bits_334;
  assign padr_bits_334 = 0;
  wire [18-1:0] padl_335;
  wire [17-1:0] padl_bits_336;
  wire [101-1:0] truncR_337;
  wire [174-1:0] truncval_338;
  wire [174-1:0] padl_339;
  wire [97-1:0] padl_bits_340;
  wire [97-1:0] padl_341;
  wire [60-1:0] padl_bits_342;
  wire [1-1:0] toSInt_343;
  assign toSInt_343 = 0;
  wire [60-1:0] toSInt_imm_344;
  wire [59-1:0] const_345;
  assign const_345 = 57646075;
  assign toSInt_imm_344 = { toSInt_343, const_345 };
  assign padl_bits_342 = toSInt_imm_344;
  assign padl_341 = { { 37{ padl_bits_342[59] } }, padl_bits_342 };
  assign padl_bits_340 = padl_341;
  assign padl_339 = { { 77{ padl_bits_340[96] } }, padl_bits_340 };
  wire [174-1:0] padl_346;
  wire [97-1:0] padl_bits_347;
  wire [97-1:0] padr_348;
  wire [59-1:0] padr_bits_349;
  assign padr_bits_349 = 0;
  assign padr_348 = { dodt, padr_bits_349 };
  assign padl_bits_347 = padr_348;
  assign padl_346 = { { 77{ padl_bits_347[96] } }, padl_bits_347 };
  assign truncval_338 = padl_339 * padl_346;
  wire [101-1:0] truncval_imm_350;
  assign truncval_imm_350 = { truncval_338[173], truncval_338[99:0] };
  assign truncR_337 = truncval_imm_350;
  wire [17-1:0] truncR_shift_351;
  assign truncR_shift_351 = truncR_337 >>> 84;
  wire [17-1:0] truncR_imm_352;
  assign truncR_imm_352 = (truncR_337[100])? truncR_shift_351[16:0] : truncR_337[100:84];
  assign padl_bits_336 = truncR_imm_352;
  assign padl_335 = { { 1{ padl_bits_336[16] } }, padl_bits_336 };
  assign padr_333 = { padl_335, padr_bits_334 };
  assign padr_331 = { padr_333, padr_bits_332 };
  assign truncval_330 = padr_331;
  wire [39-1:0] truncval_imm_353;
  assign truncval_imm_353 = { truncval_330[40], truncval_330[37:0] };

  always @(posedge clk) begin
    prev_sys_clk <= sys_clk;
  end

  localparam fsm_1 = 1;
  localparam fsm_2 = 2;
  localparam fsm_3 = 3;
  localparam fsm_4 = 4;

  always @(posedge clk) begin
    if(reset) begin
      fsm <= fsm_init;
    end else begin
      case(fsm)
        fsm_init: begin
          if(reset) begin
            o <= 39'd226774273228;
          end else begin
            o <= padr_0;
          end
          if(~prev_sys_clk & sys_clk & ((VREF > VREG) & (VREF <= 15'd16384))) begin
            fsm <= fsm_1;
          end 
        end
        fsm_1: begin
          if(reset) begin
            o <= 39'd226774273228;
          end else begin
            o <= padr_57;
          end
          if(state_cycle_counter > wait_time) begin
            state_cycle_counter <= 0;
          end else begin
            state_cycle_counter <= state_cycle_counter + 1;
          end
          if(state_cycle_counter > wait_time) begin
            fsm <= fsm_2;
          end 
        end
        fsm_2: begin
          if(reset) begin
            o <= 39'd226774273228;
          end else begin
            o <= o + truncval_imm_173;
          end
          if(prev_sys_clk & ~sys_clk) begin
            fsm <= fsm_3;
          end 
        end
        fsm_3: begin
          if(reset) begin
            o <= 39'd226774273228;
          end else begin
            o <= padl_231;
          end
          if(state_cycle_counter > wait_time_lh) begin
            state_cycle_counter <= 0;
          end else begin
            state_cycle_counter <= state_cycle_counter + 1;
          end
          if(state_cycle_counter > wait_time_lh) begin
            fsm <= fsm_4;
          end 
        end
        fsm_4: begin
          if(reset) begin
            o <= 39'd226774273228;
          end else begin
            o <= o + truncval_imm_353;
          end
          if((o > 39'd226087078461) & (o <= 39'd274877906944)) begin
            fsm <= fsm_init;
          end 
        end
      endcase
    end
  end


endmodule

